
//Exercicio 4 Design


module sillyfunction (
	input logic a, b,
	output logic y);

	assign y = a ^ b;
endmodule